module async_fifo_top #(
    parameter DATA_WIDTH = 8,
    parameter ADDR_WIDTH = 4
)(
    // --- Write Domain ---
    input  logic                  w_clk,
    input  logic                  w_rst_n,
    input  logic                  w_inc,
    input  logic [DATA_WIDTH-1:0] w_data,
    output logic                  w_full,

    // --- Read Domain ---
    input  logic                  r_clk,
    input  logic                  r_rst_n,
    input  logic                  r_inc,
    output logic [DATA_WIDTH-1:0] r_data,
    output logic                  r_empty
);

    logic [ADDR_WIDTH-1:0] w_addr, r_addr;
    logic [ADDR_WIDTH:0]   w_ptr, r_ptr;
    logic [ADDR_WIDTH:0]   w_q2_r_ptr, r_q2_w_ptr;

    // 1. CDC: Read -> Write (sync_2ff yerine multi_ff kullanıyoruz)
    multi_ff #(.WIDTH(ADDR_WIDTH+1)) sync_r2w (
        .clk   (w_clk),
        .rst_n (w_rst_n),
        .IN_0  (r_ptr),       // multi_ff port ismi
        .OUT_1 (w_q2_r_ptr)   // multi_ff port ismi
    );

    // 2. CDC: Write -> Read
    multi_ff #(.WIDTH(ADDR_WIDTH+1)) sync_w2r (
        .clk   (r_clk),
        .rst_n (r_rst_n),
        .IN_0  (w_ptr),       // multi_ff port ismi
        .OUT_1 (r_q2_w_ptr)   // multi_ff port ismi
    );

    // 3. Write Logic
    w_ptr_full_flag #(.ADDR_WIDTH(ADDR_WIDTH)) w_ptr_handler (
        .w_clk      (w_clk),
        .w_rst_n    (w_rst_n),
        .w_inc      (w_inc),
        .w_q2_r_ptr (w_q2_r_ptr),
        .w_full     (w_full),
        .w_addr     (w_addr),
        .w_ptr      (w_ptr)
    );

    // 4. Read Logic
    r_ptr_empty_flag #(.ADDR_WIDTH(ADDR_WIDTH)) r_ptr_handler (
        .r_clk      (r_clk),
        .r_rst_n    (r_rst_n),
        .r_inc      (r_inc),
        .r_q2_w_ptr (r_q2_w_ptr),
        .r_empty    (r_empty),
        .r_addr     (r_addr),
        .r_ptr      (r_ptr)
    );

    // 5. Memory
    mem #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH)
    ) fifo_ram (
        .w_clk   (w_clk),
        .w_inc   (w_inc),
        .w_full  (w_full),
        .w_addr  (w_addr),
        .w_data  (w_data),
        
        .r_clk   (r_clk),
        .r_inc   (r_inc),
        .r_empty (r_empty),
        .r_addr  (r_addr),
        .r_data  (r_data)
    );

endmodule